library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity sinerom is
    Port ( addr : in std_logic_vector(7 downto 0);
           sin : out std_logic_vector(7 downto 0));
end sinerom;

architecture Behavioral of sinerom is

type SINROM is array (0 to 255) of STD_LOGIC_VECTOR(7 downto 0);

constant ROMVALS : SINROM := ("10000000","10000011","10000110","10001001",
                              "10001100","10010000","10010011","10010110",
                              "10011001","10011100","10011111","10100010",
						"10100101","10101000","10101011","10101110",
						"10110001","10110011","10110110","10111001",
						"10111100","10111110","11000001","11000100",
						"11000110","11001001","11001100","11001110",
						"11010000","11010011","11010101","11010111",
						"11011010","11011100","11011110","11100000",
						"11100010","11100100","11100110","11101000",
						"11101001","11101011","11101101","11101110",
						"11110000","11110001","11110011","11110100",
						"11110101","11110110","11110111","11111001",
						"11111001","11111010","11111011","11111100",
						"11111100","11111101","11111110","11111110",
						"11111110","11111111","11111111","11111111",
						"11111111","11111111","11111111","11111111",
						"11111110","11111110","11111110","11111101",
						"11111101","11111100","11111011","11111011",
						"11111010","11111001","11111000","11110111",
						"11110110","11110100","11110011","11110010",
						"11110000","11101111","11101101","11101100",
						"11101010","11101000","11100110","11100100",
						"11100010","11100001","11011110","11011100",
						"11011010","11011000","11010110","11010011",
						"11010001","11001111","11001100","11001010",
						"11000111","11000100","11000010","11000000",
						"10111100","10111010","10110111","10110100",
						"10110001","10101110","10101011","10101000",
						"10100101","10100010","10011111","10011100",
						"10011001","10010110","10010011","10010000",
						"10001101","10001010","10000111","10000100",
						"10000001","10000000","01111010","01110111",
						"01110100","01110001","01101110","01101011",
						"01101000","01100101","01100010","01011111",
						"01011100","01011001","01010110","01010011",
						"01010000","01001101","01001010","01001000",
						"01000101","01000010","00111111","00111101",
						"00111010","00111000","00110101","00110011",
						"00110000","00101110","00101011","00101001",
						"00100111","00100101","00100011","00100000",
						"00011110","00011100","00011011","00011001",
						"00010111","00010101","00010100","00010010",
						"00010000","00001111","00001110","00001100",
						"00001011","00001010","00001001","00001000",
						"00000111","00000110","00000101","00000100",
						"00000100","00000011","00000011","00000010",
						"00000010","00000001","00000001","00000001",
						"00000001","00000001","00000001","00000001",
						"00000010","00000010","00000010","00000011",
						"00000011","00000100","00000101","00000101",
						"00000110","00000111","00001000","00001001",
						"00001010","00001011","00001101","00001110",
						"00001111","00010001","00010010","00010100",
						"00010110","00010111","00011001","00011011",
						"00011101","00011111","00100001","00100011",
						"00100101","00101000","00101010","00101100",
						"00101110","00110001","00110011","00110110",
						"00111000","00111011","00111110","01000000",
						"01000011","01000110","01001001","01001011",
						"01001110","01010001","01010100","01010111",
						"01011010","01011101","01100000","01100011",
						"01100110","01101001","01101100","01101111",
						"01110010","01110101","01111000","01111011");
begin
  sin <= ROMVALS(conv_integer(addr));
end Behavioral;